`timescale 1ns / 1ps

module tb_d_ff();
    reg din,clk,rst;
    wire dout;
    
    
    
    
endmodule
